//`ifndef __RSA__DEFINE__
//`define __RSA__DEFINE__
// 128, 256, 512, 1024
parameter RSA_BIT_MAX = 11'd1024;
parameter RSA_BIT_LOG2_MAX = 4'd10;
//`endif