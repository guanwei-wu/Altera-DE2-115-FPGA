//`ifndef __RSA__DEFINE__
//`define __RSA__DEFINE__
// 128, 256, 512, 1024
parameter RSA_BIT_MAX = 10'd512;
parameter RSA_BIT_LOG2_MAX = 4'd9;
//`endif